//
// File Name: alucodes.sv
// Function: ALU codes
// Author: Mohammad Abu Alhalawe
// Last rev.: 05/09/19
//
`define	alu_add   5'h00
`define	alu_addu  5'h01
`define	alu_sltu  5'h02
`define	alu_subu  5'h03
`define	alu_slli  5'h04
`define	alu_srli  5'h05
`define	alu_srai  5'h06
`define	alu_sub   5'h07
`define	alu_and   5'h08
`define	alu_or    5'h09
`define	alu_xor   5'h0A
`define	alu_sll   5'h0B
`define	alu_srl   5'h0C
`define	alu_sra   5'h0D
`define	alu_nor   5'h0E
`define  alu_slt  5'h0F
`define alu_mul   5'h10
`define alu_div   5'h11
`define alu_mulh  5'h12
`define alu_divu  5'h13
`define alu_rem   5'h14
`define alu_remu  5'h15
`define alu_mulhu 5'h16
