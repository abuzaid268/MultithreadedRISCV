@0
0000000A
00000009
00000008 
00000007 
00000006
00000005 
00000004 
00000003 
00000002 
00000001 
00000001 
00000002 
00000003 
00000004 
00000005 
00000006 
00000007 
00000008 
00000009 
0000000A 
00000009
00000008
00000007
00000006
00000005
00000004
00000003
00000002
00000001
00000000
00000000
00000001
00000002
00000003
00000004
00000005
00000006
00000007
00000008
00000009
00000009
00000008
00000007
00000006
00000005
00000004
00000003
00000002
00000001
00000000