@00000000
73 62 40 F1 93 02 00 00 13 03 10 00 93 03 20 00 
13 0E 30 00 63 04 52 00 6F 00 40 01 37 21 00 00 
37 24 00 00 93 00 00 00 6F 00 00 04 63 04 62 00 
6F 00 40 01 37 41 00 00 37 44 00 00 93 00 00 00 
6F 00 80 02 63 04 72 00 6F 00 40 01 37 61 00 00 
37 64 00 00 93 00 00 00 6F 00 00 01 37 81 00 00 
37 84 00 00 93 00 00 00 13 01 01 FD 23 26 11 02 
23 24 81 02 13 04 01 03 23 22 04 FE 23 20 04 FE 
23 2E 04 FC 23 2C 04 FC 23 2A 04 FE 23 28 04 FE 
23 26 04 FE 23 24 04 FE F3 67 40 F1 23 2A F4 FC 
83 27 44 FD 63 9C 07 02 03 25 44 FF EF 00 80 10 
23 22 A4 FE 13 07 00 00 83 27 44 FE 23 20 F7 00 
93 07 20 00 03 27 44 FF 23 A0 E7 00 83 27 44 FF 
93 87 17 00 23 2A F4 FE 6F F0 1F FD 03 27 44 FD 
93 07 10 00 63 1C F7 02 03 25 04 FF EF 00 80 11 
23 20 A4 FE 93 07 40 00 03 27 04 FE 23 A0 E7 00 
93 07 60 00 03 27 04 FF 23 A0 E7 00 83 27 04 FF 
93 87 17 00 23 28 F4 FE 6F F0 1F FD 03 27 44 FD 
93 07 20 00 63 1C F7 02 03 25 C4 FE EF 00 00 15 
23 2E A4 FC 93 07 80 00 03 27 C4 FD 23 A0 E7 00 
93 07 A0 00 03 27 C4 FE 23 A0 E7 00 83 27 C4 FE 
93 87 17 00 23 26 F4 FE 6F F0 1F FD 03 27 44 FD 
93 07 30 00 63 1C F7 02 03 25 84 FE EF 00 00 16 
23 2C A4 FC 93 07 C0 00 03 27 84 FD 23 A0 E7 00 
93 07 E0 00 03 27 84 FE 23 A0 E7 00 83 27 84 FE 
93 87 17 00 23 24 F4 FE 6F F0 1F FD 93 07 00 00 
13 85 07 00 83 20 C1 02 03 24 81 02 13 01 01 03 
67 80 00 00 13 01 01 FF 23 26 11 00 23 24 81 00 
13 04 01 01 23 2A A4 FE 83 27 44 FF 63 96 07 00 
93 07 00 00 6F 00 C0 01 83 27 44 FF 93 87 F7 FF 
13 85 07 00 EF F0 1F FD 93 07 05 00 93 87 37 00 
13 85 07 00 83 20 C1 00 03 24 81 00 13 01 01 01 
67 80 00 00 13 01 81 FE 23 2A 11 00 23 28 81 00 
23 26 91 00 13 04 81 01 23 26 A4 FE 83 27 C4 FE 
63 88 07 00 03 27 C4 FE 93 07 10 00 63 16 F7 00 
83 27 C4 FE 6F 00 00 03 83 27 C4 FE 93 87 F7 FF 
13 85 07 00 EF F0 1F FC 93 04 05 00 83 27 C4 FE 
93 87 E7 FF 13 85 07 00 EF F0 DF FA 93 07 05 00 
B3 87 F4 00 13 85 07 00 83 20 41 01 03 24 01 01 
83 24 C1 00 13 01 81 01 67 80 00 00 13 01 01 FF 
23 26 11 00 23 24 81 00 13 04 01 01 23 2A A4 FE 
83 27 44 FF 63 96 07 00 93 07 00 00 6F 00 C0 01 
83 27 44 FF 93 87 F7 FF 13 85 07 00 EF F0 1F FD 
93 07 05 00 93 87 47 00 13 85 07 00 83 20 C1 00 
03 24 81 00 13 01 01 01 67 80 00 00 13 01 01 FF 
23 26 11 00 23 24 81 00 13 04 01 01 23 2A A4 FE 
83 27 44 FF 63 96 07 00 93 07 00 00 6F 00 00 02 
83 27 44 FF 93 87 F7 FF 13 85 07 00 EF F0 1F FD 
13 07 05 00 83 27 44 FF B3 07 F7 00 13 85 07 00 
83 20 C1 00 03 24 81 00 13 01 01 01 67 80 00 00 
