//
// File Name: opcode.sv
// Function: instruction opcode
// Author: Mohammad Abu Alhalawe
// Last rev.: 05/09/19
//
`define LUI    7'b0110111 
`define AUIPC  7'b0010111 
`define JAL     7'b1101111
`define JALR    7'b1100111
`define Btype   7'b1100011
`define LW       7'b0000011
`define SW       7'b0100011
`define Itype    7'b0010011
`define Rtype    7'b0110011
`define Enquiry  7'b1111111
`define CSRRS    7'b1110011

